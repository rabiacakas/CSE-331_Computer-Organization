library verilog;
use verilog.vl_types.all;
entity likeALU_testbench is
end likeALU_testbench;
