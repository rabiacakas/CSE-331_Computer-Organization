library verilog;
use verilog.vl_types.all;
entity mips_core_testbench is
end mips_core_testbench;
