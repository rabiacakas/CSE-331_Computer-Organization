library verilog;
use verilog.vl_types.all;
entity mips_registers_testbench is
end mips_registers_testbench;
