library verilog;
use verilog.vl_types.all;
entity ALU_testbench is
end ALU_testbench;
